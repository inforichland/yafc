library IEEE;
use IEEE.STD_LOGIC_1164.all;

package uart_pkg is

  -- Data types
  type uart_in_ctrl is record
  end record;
  
  type uart_out_ctrl is record
  end record;

end uart_pkg;

package body uart_pkg is
end uart_pkg;
